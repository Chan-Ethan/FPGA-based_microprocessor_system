`ifndef GLOBAL_EVENTS_PKG_SVH
`define GLOBAL_EVENTS_PKG_SVH

package global_events_pkg;
  event reset_e;        // Mouse master reset command event
  event start_stream_e; // Mouse master start stream command event
endpackage

`endif // GLOBAL_EVENTS_PKG_SVH
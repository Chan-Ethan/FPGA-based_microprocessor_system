module MouseMasterSM(
input CLK,
input RESET,

//Transmitter Control
output reg          SEND_BYTE,
output reg  [7:0]   BYTE_TO_SEND,
input               BYTE_SENT,

//Receiver Control
output reg          READ_ENABLE,
input       [7:0]   BYTE_READ,
input       [1:0]   BYTE_ERROR_CODE,
input               BYTE_READY,

//Data Registers
output reg  [7:0]   MOUSE_DX,
output reg  [7:0]   MOUSE_DY,
output reg  [7:0]   MOUSE_STATUS,

output reg          SEND_INTERRUPT,
input               INTERRUPT_ACK,

// Debug signals
output      [6:0]   current_state
);

`define FSM_IDLE            7'b0000001
`define FSM_RESET           7'b0000010
`define FSM_WAIT_ACK        7'b0000100
`define FSM_WAIT_SELFTST    7'b0001000
`define FSM_STAR_STM        7'b0010000
`define FSM_WAIT_ACK2       7'b0100000
`define FSM_STREAM_MOD      7'b1000000

`ifdef SIMULATION
    `define CNT_NUM_10MS    20'd99_999
`else
    `define CNT_NUM_10MS    20'd999_999
`endif

`define CNT_BYTES       2'b10

logic [6:0]         current_state, next_state;
logic               waiting_wr_done;
logic [1:0]         byte_cnt;
logic [19:0]        cnt_10ms;
logic [23:0]        pkt_buffer;

// State Transition Logic
always_comb begin
    next_state = current_state;
    case (current_state)
        `FSM_IDLE: begin
            // Wait for the first byte to be sent and mouse initialization
            if (cnt_10ms == `CNT_NUM_10MS) next_state = `FSM_RESET;
        end
        `FSM_RESET: begin
            // send reset command
            if (BYTE_SENT) next_state = `FSM_WAIT_ACK;
        end
        `FSM_WAIT_ACK: begin
            // wait for the ack from mouse
            if (BYTE_READY) begin
                if (BYTE_ERROR_CODE != 2'b00) begin
                    next_state = `FSM_RESET;
                end
                else if (BYTE_READ == 8'hFA || BYTE_READ == 8'hF4) begin
                    next_state = `FSM_WAIT_SELFTST;
                end
                else begin
                    next_state = `FSM_RESET;
                end
            end
            else if (cnt_10ms == `CNT_NUM_10MS) begin
                next_state = `FSM_RESET;
            end
        end
        `FSM_WAIT_SELFTST: begin
            // wait for the self test packet from mouse
            if (BYTE_READY) begin
                if (BYTE_ERROR_CODE != 2'b00) begin
                    next_state = `FSM_RESET;
                end
                else if (BYTE_READ == 8'hAA) begin
                    next_state = `FSM_STAR_STM;
                end
                else begin
                    next_state = `FSM_RESET;
                end
            end
            else;
        end
        `FSM_STAR_STM: begin
            // send start streaming mode command
            if (BYTE_SENT) next_state = `FSM_WAIT_ACK2;
        end
        `FSM_WAIT_ACK2: begin
            // wait for the ack from mouse
            if (BYTE_READY) begin
                if (BYTE_ERROR_CODE != 2'b00) begin
                    next_state = `FSM_RESET;
                end
                else if (BYTE_READ == 8'hFA || BYTE_READ == 8'hF4) begin
                    next_state = `FSM_STREAM_MOD;
                end
                else begin
                    next_state = `FSM_RESET;
                end
            end
        end
        `FSM_STREAM_MOD: begin
            // keep receiving data from mouse
            if ((BYTE_READY == 1'b1) && (BYTE_ERROR_CODE != 2'b00)) begin
                // if error packet received, reset
                next_state = `FSM_RESET;
            end
            else;
        end
        default: next_state = `FSM_RESET;
    endcase
end

// State Register
always_ff @(posedge CLK or negedge RESET) begin
    if (!RESET) current_state <= `FSM_IDLE;
    else current_state <= next_state;
end

//================= Counters =================//
always_ff @(posedge CLK or negedge RESET) begin
    if (!RESET) begin
        cnt_10ms <= 20'd0;
    end
    else begin
        cnt_10ms <= (cnt_10ms == `CNT_NUM_10MS) ? 20'd0 : cnt_10ms + 20'd1;
    end
end

//================= Transmitter Control =================//
always_ff @(posedge CLK or negedge RESET) begin
    if (!RESET) begin
        SEND_BYTE <= 1'b0;
        waiting_wr_done <= 1'b0;
    end else begin
        if ((current_state == `FSM_STAR_STM) || (current_state == `FSM_RESET)) begin
            SEND_BYTE <= ~waiting_wr_done;
            waiting_wr_done <= 1'b1;
        end else begin
            SEND_BYTE <= 1'b0;
            waiting_wr_done <= 1'b0;
        end
    end
end

always@(posedge CLK or negedge RESET) begin
    if (!RESET) begin
        BYTE_TO_SEND <= 8'hFF;
    end
    else begin
        BYTE_TO_SEND <= (current_state == `FSM_STAR_STM) ? 8'hF4 : 8'hFF;
    end
end 

//================= Receiver Control =================//
always @(posedge CLK or negedge RESET) begin
    if (!RESET) begin
        READ_ENABLE <= 1'b0;
    end
    else begin
        READ_ENABLE <= (current_state != `FSM_RESET) && (current_state != `FSM_STAR_STM);
    end
end 

//================= Data Packing =================//
always_ff @(posedge CLK or negedge RESET) begin
    if (!RESET) begin
        pkt_buffer <= 24'b0;
    end
    else if (current_state == `FSM_STREAM_MOD) begin
        if (BYTE_READY == 1'b1) begin
            case (byte_cnt)
                2'b00: pkt_buffer[7:0] <= BYTE_READ;
                2'b01: pkt_buffer[15:8] <= BYTE_READ;
                2'b10: pkt_buffer[23:16] <= BYTE_READ;
                default: ;
            endcase
        end
        else;
    end
    else begin
        pkt_buffer <= 24'b0;
    end
end

always @(posedge CLK or negedge RESET) begin
    if (!RESET) begin
        byte_cnt <= 2'b00;
    end
    else if (current_state == `FSM_STREAM_MOD) begin
        if (BYTE_READY == 1'b1) begin
            byte_cnt <= (byte_cnt == `CNT_BYTES) ? 2'b00 : byte_cnt + 2'b01;
        end
        else;
    end
    else begin
        byte_cnt <= 2'b00;
    end

end


//================= Output Registers =================//
assign MOUSE_STATUS = pkt_buffer[7:0];
assign MOUSE_DX = pkt_buffer[15:8];
assign MOUSE_DY = pkt_buffer[23:16];

always @(posedge CLK or negedge RESET) begin
    if (!RESET) begin
        SEND_INTERRUPT <= 1'b0;
    end
    else if (INTERRUPT_ACK == 1'b1) begin
        SEND_INTERRUPT <= 1'b0;
    end
    else if ((current_state == `FSM_STREAM_MOD) && 
             (BYTE_READY == 1'b1) && 
             (byte_cnt == `CNT_BYTES)) begin
        SEND_INTERRUPT <= 1'b1;
    end
    else;
end

endmodule
